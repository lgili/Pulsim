* RL Step Response - LTspice benchmark
* Matches Pulsim benchmarks/circuits/rl_step.yaml

V1 in 0 PULSE(0 10 0 1n 1n 10m 20m)
R1 in out 100
L1 out 0 10m IC=0

.tran 1u 1m UIC
.backanno
.end
