* RC Low-pass Filter - LTspice benchmark
* Matches Pulsim benchmarks/circuits/rc_dc.yaml

V1 in 0 DC 5.0
R1 in out 1k
C1 out 0 1u IC=0

.tran 1u 5m UIC
.backanno
.end
